/* Verilog model created from schematic sch_test.sch -- Oct 19, 2013 21:09 */

module sch_test;




endmodule // sch_test
